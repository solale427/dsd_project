`timescale 1ns / 1ps

module tbt_fbf_adder_tb();
    reg A_stb_tbt;
    reg B_stb_tbt;
    reg clk;
    reg reset;
    reg result_ack_tbt;
    reg [32 * 2 * 2 - 1:0] A_tbt;
    reg [32 * 2 * 2 - 1:0] B_tbt;
    wire result_ready_tbt;
    wire [32 * 2 * 2 - 1:0] result_tbt;
    
    reg A_stb_fbf;
    reg B_stb_fbf;
    reg result_ack_fbf;
    reg [32 * 4 * 4 - 1:0] A_fbf;
    reg [32 * 4 * 4 - 1:0] B_fbf;
    wire result_ready_fbf;
    wire [32 * 4 * 4 - 1:0] result_fbf;
    reg [31:0] result_tbt_2d_array[1:0][1:0];
    reg [127:0] correct_result_tbt;
    reg [511:0] correct_result_fbf;
    
    tbt_adder tbtAdder (
    .A_stb(A_stb_tbt),
    .B_stb(B_stb_tbt),
    .clk(clk),
    .reset(reset),
    .result_ack(result_ack_tbt),
    .A(A_tbt),
    .B(B_tbt),
    .result_ready(result_ready_tbt),
    .result(result_tbt)
);
    fbf_adder fbfAdder (
    .A_stb(A_stb_fbf),
    .B_stb(B_stb_fbf),
    .clk(clk),
    .reset(reset),
    .result_ack(result_ack_fbf),
    .A(A_fbf),
    .B(B_fbf),
    .result_ready(result_ready_fbf),
    .result(result_fbf)
);

    initial
   begin
      clk = 0;
      forever
        #10 clk = ~clk;
   end

initial begin
reset = 0;
#12;
reset = 1;
A_stb_tbt = 1;
B_stb_tbt = 1;
A_stb_fbf = 1;
B_stb_fbf = 1;
$monitor("result_ready_tbt = %b, result_ready_fbf = %b, result_tbt = %h, correct_result_tbt = %h, result_fbf = %h, correct_result_fbf = %h ",
            result_ready_tbt,
            result_ready_fbf,
            result_tbt,
            correct_result_tbt,
            result_fbf,
            correct_result_fbf
            );
            
    //	A_mtrix_form = | 5.84   8.16 |
	//		           | -3.01  -10  |
	//
	//	B_matrix_form = | 20.9   -12.8|
	//		            | 9.35   2    |
	//	
	//	result_matrix_form = | 26.74  -4.64|
	//		                 | 6.34  -8|
	
    A_tbt[31:0] = 32'b01000000101110101110000101001000;
    A_tbt[63:32] = 32'b01000001000000101000111101011100; 
    A_tbt[95:64] = 32'b11000000010000001010001111010111;
    A_tbt[127:96] = 32'b11000001001000000000000000000000;
    
    B_tbt[31:0] = 32'b01000001101001110011001100110011;
    B_tbt[63:32] = 32'b11000001010011001100110011001101; 
    B_tbt[95:64] = 32'b01000001000101011001100110011010;
    B_tbt[127:96] = 32'b01000000000000000000000000000000;
    
    correct_result_tbt[31:0] = 32'b01000001110101011110101110000101;
    correct_result_tbt[63:32] = 32'b11000000100101000111101011100001;
    correct_result_tbt[95:64] = 32'b01000000110010101110000101001000;
    correct_result_tbt[127:96] = 32'b11000001000000000000000000000000;
    
    
    //	A_mtrix_form = |1.2   4.34  8.16  3.21|
	//		           |-1.9  2.3  -11  -1.5|
	//                 |-3.01  -10  21.54  -5.6|
	//                 |1.2  0.72  32  -0.98|
	//	B_matrix_form = |13.63   -12.8  11.2  1.3|
	//		            |8.35   2  4.3  6.78|
	//		            |-4.1   -8.76   8.16  -9.75 |
	//		            |-2.12  6.34  1.98  13.4 |

	//	result_matrix_form = |14.83  -8.46  19.36  4.51|
	//		                 |6.45  4.3  -6.7  5.28|
	//		                 |-7.11  -18.76  29.7  15.35|
	//		                 |-0.92  7.06  33.98  12.42|
		   
    A_fbf[31:0] = 32'b00111111100110011001100110011010;
    A_fbf[63:32] = 32'b01000000100010101110000101001000; 
    A_fbf[95:64] = 32'b01000001000000101000111101011100;
    A_fbf[127:96] = 32'b01000000010011010111000010100100;
    A_fbf[159:128] = 32'b10111111111100110011001100110011;
    A_fbf[191:160] = 32'b01000000000100110011001100110011;
    A_fbf[223:192] = 32'b11000001001100000000000000000000;
    A_fbf[255:224] = 32'b10111111110000000000000000000000;
    A_fbf[287:256] = 32'b11000000010000001010001111010111;
    A_fbf[319:288] = 32'b11000001001000000000000000000000;
    A_fbf[351:320] = 32'b01000001101011000101000111101100;
    A_fbf[383:352] = 32'b11000000101100110011001100110011;
    A_fbf[415:384] = 32'b00111111100110011001100110011010;
    A_fbf[447:416] = 32'b00111111001110000101000111101100;
    A_fbf[479:448] = 32'b01000010000000000000000000000000;
    A_fbf[511:480] = 32'b10111111011110101110000101001000;
    
    B_fbf[31:0] = 32'b01000001010110100001010001111011;
    B_fbf[63:32] = 32'b11000001010011001100110011001101; 
    B_fbf[95:64] = 32'b01000001001100110011001100110011;
    B_fbf[127:96] = 32'b00111111101001100110011001100110;
    B_fbf[159:128] = 32'b01000001000001011001100110011010;
    B_fbf[191:160] = 32'b01000000000000000000000000000000;
    B_fbf[223:192] = 32'b01000000100010011001100110011010;
    B_fbf[255:224] = 32'b01000000110110001111010111000011;
    B_fbf[287:256] = 32'b11000000100000110011001100110011;
    B_fbf[319:288] = 32'b11000001000011000010100011110110;
    B_fbf[351:320] = 32'b01000001000000101000111101011100;
    B_fbf[383:352] = 32'b11000001000111000000000000000000;
    B_fbf[415:384] = 32'b11000000000001111010111000010100;
    B_fbf[447:416] = 32'b01000000110010101110000101001000;
    B_fbf[479:448] = 32'b00111111111111010111000010100100;
    B_fbf[511:480] = 32'b01000001010101100110011001100110;

    correct_result_fbf[31:0] = 32'b01000001011011010100011110101110;        
    correct_result_fbf[63:32] = 32'b11000001000001110101110000101001;
    correct_result_fbf[95:64] = 32'b01000001100110101110000101001000;
    correct_result_fbf[127:96] = 32'b01000000100100000101000111101100;
    correct_result_fbf[159:128] = 32'b01000000110011100110011001100110;
    correct_result_fbf[191:160] = 32'b01000000100010011001100110011010;
    correct_result_fbf[223:192] = 32'b11000000110101100110011001100110;
    correct_result_fbf[255:224] = 32'b01000000101010001111010111000011;
    correct_result_fbf[287:256] = 32'b11000000111000111000010100011111;
    correct_result_fbf[319:288] = 32'b11000001100101100001010001111011;
    correct_result_fbf[351:320] = 32'b01000001111011011001100110011010;
    correct_result_fbf[383:352] = 32'b01000001011101011001100110011010;
    correct_result_fbf[415:384] = 32'b10111111011010111000010100011111;
    correct_result_fbf[447:416] = 32'b01000000111000011110101110000101;
    correct_result_fbf[479:448] = 32'b01000010000001111110101110000101;
    correct_result_fbf[511:480] = 32'b01000001010001101011100001010010;
    
    
end
endmodule
