module fbf_multiplier_TB();

    reg clock = 0;
    reg A_stb, B_stb;
    reg reset = 1;
    reg result_ack = 0;
    reg [32 * 4 * 4 - 1:0] A, B;
	wire [3:0] state;
    wire [32 * 4 * 4 - 1:0] result;
    wire ready;
    
    initial
    begin
        forever
            #10 clock = ~clock;
    end
    
    initial
    begin
        A = 512'b01000000100010011001100110011010001111111100110011001100110011010011111011001100110011001100110100111110100110011001100110011010001111100100110011001100110011010100000011101001100110011001101001000000101110011001100110011010010000001010011001100110011001100100000011001001100110011001101001000000001000000000000000000000010000001001011001100110011001100100000000000110011001100110011001000000101010011001100110011010001111101100110011001100110011010100000000010011001100110011001100111111110000000000000000000000;
        B = 512'b01000000001000000000000000000000010000001101110011001100110011010100000000111001100110011001101001000000100011001100110011001101010000000111100110011001100110100100000010110011001100110011001101000001000111100110011001100110010000000101001100110011001100110100000011110110011001100110011001000000101000110011001100110011001111111010011001100110011001100011111111001100110011001100110101000000000001100110011001100110001111111111001100110011001100110011111111011001100110011001101000111111100011001100110011001101;
       	//A = 512'b0;
        //B = 512'b0;
        A_stb = 1;
        B_stb = 1;
        $monitor("ready: %b result: %b", ready, result);
    end
    
    fbf_multiplier multiplier(
    .A_stb(A_stb),
    .B_stb(B_stb),
    .clk(clock),
    .reset(reset),
    .result_ack(result_ack),
    .A(A),
    .B(B),
    .result_ready(ready),
    .result(result)
);

endmodule