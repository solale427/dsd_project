module sync_ram #(
  parameter ADDR_WIDTH=16             //width of addresse bus
)(
  input  [31:0] 	    Din,     //data to be written
  input  [(ADDR_WIDTH-1):0] addr,    //address for write/read operation
  input                     writeEn, //write enable signal
  input			    read,    //read enable signal
  input                     clk,     //clock signal
  output  [31:0]            Dout     //read data
);
  localparam RAM_DEPTH = 1 << ADDR_WIDTH;
  reg [31:0] mem [RAM_DEPTH-1:0];
  
  reg [42*32-1:0] A;
  reg [30*32-1:0] B;
  integer i;
  
  initial
  begin
  
    mem[0] = {31'b0, 1'b1};
    mem[1] = {8'd5, 8'd6, 8'd6, 8'd7};
    /*mem[17] = 32'b01000000100010011001100110011010;
    mem[16] = 32'b00111111110011001100110011001101;
    mem[15] = 32'b00111110110011001100110011001101;
    mem[14] = 32'b00111110100110011001100110011010;
    mem[13] = 32'b00111110010011001100110011001101;
    mem[12] = 32'b01000000111010011001100110011010;
    mem[11] = 32'b01000000101110011001100110011010;
    mem[10] = 32'b01000000101001100110011001100110;
    mem[9] = 32'b01000000110010011001100110011010;
    mem[8] = 32'b01000000001000000000000000000000;
    mem[7] = 32'b01000000100101100110011001100110;
    mem[6] = 32'b01000000000001100110011001100110;
    mem[5] = 32'b01000000101010011001100110011010;
    mem[4] = 32'b00111110110011001100110011001101;
    mem[3] = 32'b01000000000100110011001100110011;
    mem[2] = 32'b00111111110000000000000000000000;
    
    mem[10002] = 32'b00111111100011001100110011001101;
    mem[10003] = 32'b00111111110110011001100110011010;
    mem[10004] = 32'b00111111111100110011001100110011;
    mem[10005] = 32'b01000000000001100110011001100110;
    mem[10006] = 32'b00111111110011001100110011001101;
    mem[10007] = 32'b00111111101001100110011001100110;
    mem[10008] = 32'b01000000101000110011001100110011;
    mem[10009] = 32'b01000000111101100110011001100110;
    mem[10010] = 32'b01000000010100110011001100110011;
    mem[10011] = 32'b01000001000111100110011001100110;
    mem[10012] = 32'b01000000101100110011001100110011;
    mem[10013] = 32'b01000000011110011001100110011010;
    mem[10014] = 32'b01000000100011001100110011001101;
    mem[10015] = 32'b01000000001110011001100110011010;
    mem[10016] = 32'b01000000110111001100110011001101;
    mem[10017] = 32'b01000000001000000000000000000000;*/
    
    
    /*mem[2] = 32'b00111111100011001100110011001101;
    mem[3] = 32'b00111111110110011001100110011010;
    mem[4] = 32'b00111111111100110011001100110011;
    mem[5] = 32'b01000000000001100110011001100110;
    mem[6] = 32'b01000000010100110011001100110011;
    mem[7] = 32'b01000000100100000000000000000000;
    mem[8] = 32'b01000000001110011001100110011010;

    mem[9] = 32'b00111111110011001100110011001101;
    mem[10] = 32'b00111111101001100110011001100110;
    mem[11] = 32'b01000000101000110011001100110011;
    mem[12] = 32'b01000000111101100110011001100110;
    mem[13] = 32'b00111111101100110011001100110011;
    mem[14] = 32'b01000000011000000000000000000000;
    mem[15] = 32'b01000000001001100110011001100110;

    mem[16] = 32'b01000000010100110011001100110011;
    mem[17] = 32'b01000001000111100110011001100110;
    mem[18] = 32'b01000000101100110011001100110011;
    mem[19] = 32'b01000000011110011001100110011010;
    mem[20] = 32'b01000000100100000000000000000000;
    mem[21] = 32'b01000000111100110011001100110011;
    mem[22] = 32'b01000000100110011001100110011010;

    mem[23] = 32'b01000000100011001100110011001101;
    mem[24] = 32'b01000000001110011001100110011010;
    mem[25] = 32'b01000000110111001100110011001101;
    mem[26] = 32'b01000000001000000000000000000000;
    mem[27] = 32'b00111111110000000000000000000000;
    mem[28] = 32'b01000000010100110011001100110011;
    mem[29] = 32'b01000000000110011001100110011010;
    
    
    
    mem[10002] = 32'b00111111110000000000000000000000;
    mem[10003] = 32'b01000000000100110011001100110011;
    mem[10004] = 32'b00111110110011001100110011001101;
    mem[10005] = 32'b01000000101010011001100110011010;

    mem[10006] = 32'b01000000000001100110011001100110;
    mem[10007] = 32'b01000000100101100110011001100110;
    mem[10008] = 32'b01000000001000000000000000000000;
    mem[10009] = 32'b01000000110010011001100110011010;

    mem[10010] = 32'b01000000101001100110011001100110;
    mem[10011] = 32'b01000000101110011001100110011010;
    mem[10012] = 32'b01000000111010011001100110011010;
    mem[10013] = 32'b00111110010011001100110011001101;

    mem[10014] = 32'b00111110100110011001100110011010;
    mem[10015] = 32'b00111110110011001100110011001101;
    mem[10016] = 32'b00111111110011001100110011001101;
    mem[10017] = 32'b01000000100010011001100110011010;

    mem[10018] = 32'b01000000011100110011001100110011;
    mem[10019] = 32'b01000001000101100110011001100110;
    mem[10020] = 32'b01000000001011001100110011001101;
    mem[10021] = 32'b00111111110110011001100110011010;
 
    mem[10022] = 32'b01000000001000000000000000000000;
    mem[10023] = 32'b01000000001001100110011001100110;
    mem[10024] = 32'b01000000010100110011001100110011;
    mem[10025] = 32'b01000000110100000000000000000000;

    mem[10026] = 32'b01000001000101001100110011001101;
    mem[10027] = 32'b01000000010110011001100110011010;
    mem[10028] = 32'b01000000001001100110011001100110;
    mem[10029] = 32'b01000000100100000000000000000000;*/
    
    //A = 3520'b1100000001010011001100110011001101000001000011001100110011001101010000010000010011001100110011010100000011100011001100110011001111000000010100110011001100110011110000010001001100110011001100111100000100011001100110011001101001000000111001100110011001100110101111101100110011001100110011010100000010110110011001100110011011000001000110000000000000000000110000000001001100110011001100111100000011100011001100110011001101000001000010000000000000000000110000001010110011001100110011010100000000100110011001100110011001000001000100011001100110011010110000000110110011001100110011011100000010110110011001100110011011000001000111001100110011001101101111111010011001100110011001101011111100011001100110011001101001000000011110011001100110011010110000001111011001100110011001101011111110011001100110011001101001000001000011100110011001100110110000000111001100110011001100111100000100001100110011001100110110111111100000000000000000000000110000010001010011001100110011010100000011000011001100110011001101000000111101100110011001100110101111110100110011001100110011010100000010110000000000000000000011000000010000000000000000000000110000001011011001100110011001100100000010111100110011001100110111000000100000110011001100110011110000000010011001100110011001100011111110001100110011001100110111000000011000000000000000000000010000001001001100110011001100111011111110100110011001100110011000111111101100110011001100110011010000010000010011001100110011011100000010010000000000000000000001000000111101100110011001100110001111111100000000000000000000001100000100000001100110011001101011000001000000000000000000000000110000001000110011001100110011010100000001111001100110011001101001000000000001100110011001100110010000001000001100110011001100110011111100000000000000000000000011000000111001100110011001100110010000001111001100110011001100111100000000010011001100110011001111000000110011001100110011001101010000010000000000000000000000001100000000000000000000000000000011000000010000000000000000000000010000001101001100110011001100111100000100010110011001100110011001000000101000000000000000000000010000010001110011001100110011010100000010011001100110011001101000111111100110011001100110011010110000001111011001100110011001101100000100000100110011001100110111000001000001001100110011001101110000001011011001100110011001101100000100001100110011001100110101000000101001100110011001100110010000010001011001100110011001101011110111001100110011001100110111000000010001100110011001100110101111111101100110011001100110100100000000000110011001100110011011000000001110011001100110011010110000001000000000000000000000001100000100001110011001100110011001000000010011001100110011001101010000001000100110011001100110101100000010001100110011001100110111000000101001100110011001100110010000010000100000000000000000000100000001011001100110011001101011000001000101100110011001100110010000001011000000000000000000001011111100110011001100110011001111000000000100110011001100110011101111110001100110011001100110100100000010110011001100110011001101000001000111001100110011001101110000001001011001100110011001101011111010011001100110011001101001000001000010000000000000000000001111111010011001100110011001100100000100011011001100110011001111000000010000000000000000000000010000010000011001100110011001100011111101100110011001100110011011000000110000000000000000000000010000010000100000000000000000001100000011110011001100110011001111000001000110000000000000000000110000010001100000000000000000001100000010010000000000000000000001000001000010000000000000000000;
    
    //B = 4160'b01000000101111001100110011001101010000000000110011001100110011011011111110001100110011001100110111000000101100000000000000000000110000010001011001100110011001101100000001001100110011001100110110111101110011001100110011001101110000001101100110011001100110101100000100011100110011001100110101000000101000110011001100110011010000010001000110011001100110101100000100000110011001100110011011000001000010000000000000000000110000001110011001100110011001101100000010001001100110011001101011000000000001100110011001100110101111110000000000000000000000000100000100011110011001100110011000111111000110011001100110011010010000001100001100110011001100110011111110110011001100110011001101000000101000110011001100110011110000001101110011001100110011011100000011001100110011001100110111000000010000000000000000000000110000000000110011001100110011011100000100001000000000000000000011000000101010011001100110011010010000000101001100110011001100110100000100010001100110011001101001000001000011001100110011001101101111110110011001100110011001101100000000011001100110011001101001000000110011001100110011001101001111111011001100110011001100111100000001000000000000000000000011000000000001100110011001100110001111100100110011001100110011010100000011110000000000000000000001000000000100110011001100110011110000001010011001100110011001101100000011100000000000000000000011000001000010000000000000000000110000001110110011001100110011010100000010000011001100110011001101000000110011001100110011001101110000001000110011001100110011011100000011100011001100110011001100111111100000000000000000000000110000010001010011001100110011010100000011000011001100110011001101000000111010011001100110011010010000001011100110011001100110101100000000000110011001100110011001000000010001100110011001100110110000000101001100110011001100110100000011010000000000000000000011000000111101100110011001100110110000001101110011001100110011010100000100000001100110011001101011000000110111001100110011001101110000001010100110011001100110100100000001110011001100110011001101000001000001100110011001100110101111111100110011001100110011011100000001010011001100110011001111000000010011001100110011001101010000000000110011001100110011011011111010011001100110011001101011000001000000110011001100110011110000001001000000000000000000001100000100000001100110011001101011000000110110011001100110011010010000001100100110011001100110101100000100011110011001100110011011000001000111100110011001100110110000001010100110011001100110100100000011011100110011001100110101000000101100000000000000000000110000001101110011001100110011010100000010101100110011001100110111000001000111100110011001100110110000001110011001100110011001101100000011010011001100110011001101000000101011001100110011001101110000010001100110011001100110100100000001010011001100110011001101000001000010000000000000000000110000001111000000000000000000001100000010100011001100110011001101000001000000000000000000000000110000010000100110011001100110101100000000110011001100110011001111000001000110000000000000000000010000000100000000000000000000001100000011110011001100110011001101000000100110011001100110011010110000010001011001100110011001100100000001000110011001100110011011000000111011001100110011001101001111110001100110011001100110100100000000000000000000000000000011000001000000110011001100110011010000010001010011001100110011010100000010100011001100110011001101000001000100011001100110011010010000010000000110011001100110100100000010100110011001100110011001000000110001100110011001100110110000000010011001100110011001101100000100011100110011001100110111000000011011001100110011001101101111110110011001100110011001101100000000000110011001100110011011000000001100110011001100110011110000001111110011001100110011010100000010100011001100110011001111000000010110011001100110011010001111111111001100110011001100111100000011010000000000000000000011000000101110011001100110011010110000001011000000000000000000000011111100000000000000000000000011000001000100000000000000000000010000001101110011001100110011010100000100001001100110011001101011000001000000011001100110011010101111111101100110011001100110100100000100000011001100110011001100111111100000000000000000000000;
    
	A = 1344'b110000010000010011001100110011011100000010010000000000000000000011000000001001100110011001100110001111111110011001100110011001100011111101001100110011001100110101000000100100110011001100110011010000000011100110011001100110101011111110100110011001100110011000111111110011001100110011001101110000010000101100110011001100111100000010110000000000000000000001000000000011001100110011001101010000001101100110011001100110100100000000001100110011001100110100111111101100110011001100110011010000000100110011001100110011010100000100011000000000000000000000111111110110011001100110011010010000001111001100110011001100110100000010100110011001100110011011000000011011001100110011001101010000001001110011001100110011010100000011010011001100110011001111000000111100110011001100110011110000001000110011001100110011011011111100011001100110011001101001000000110000110011001100110011010000010001011001100110011001101011111100011001100110011001101001000000110110011001100110011010110000001110001100110011001100111100000011000110011001100110011011000001000010000000000000000000110000001110100110011001100110101100000100000110011001100110011011000000111000000000000000000000010000010000001100110011001100110011111010011001100110011001101001000000101011001100110011001101010000001000011001100110011001100011111111011001100110011001101000111111001100110011001100110011;
	B =  960'b010000010000111001100110011001101100000100000011001100110011001100111111101100110011001100110011010000000010000000000000000000000100000011100110011001100110011001000001000101100110011001100110010000001001011001100110011001100100000010100110011001100110011001000000100000110011001100110011110000000111100110011001100110101011111011001100110011001100110111000000100011001100110011001101110000010000010011001100110011011100000001011001100110011001101010111111111001100110011001100110101111111111001100110011001100111100000011001100110011001100110111000000000000000000000000000000110000000100110011001100110011011100000001101100110011001100110101000000101100110011001100110011110000001111000000000000000000000100000010000110011001100110011001000001000010011001100110011010101111101100110011001100110011010100000010001100110011001100110111000000010011001100110011001101101111111110011001100110011001101100000001111001100110011001101001000000100000000000000000000000;	

    for(i = 0; i < 42; i = i + 1)
    begin
        mem[i + 2] = A[(1343-i*32)-:32];
    end
    
    for(i = 0; i < 30; i = i + 1)
    begin
        mem[i + 10002] = B[(959-i*32)-:32];
    end
    
  end
  
  
  
  assign Dout = (read) ? mem[addr] : 32'bz;

  always @(posedge clk) begin //WRITE
      if (writeEn) begin
          mem[addr] <= Din;
      end
  end
  
endmodule