`timescale 1ns / 1ps

module fbf_testbench
#(
	parameter FLOAT_SIZE = 32
)
();


parameter zero = 32'b00000000000000000000000000000000;
parameter one = 32'b00111111100000000000000000000000;
reg clk = 1'b0;
reg [16*FLOAT_SIZE-1:0] A;
reg [16*FLOAT_SIZE-1:0] B;
wire [16*FLOAT_SIZE-1:0] Res; 
wire ready;
reg load = 1'b0;
reg reset = 1'b1;
reg A_stb = 1'b0;
reg B_stb = 1'b0;
reg result_ack = 1'b0;

fbf_multiplier fbf_mult_test(
	.clk(clk),
	.reset(reset),
	.A(A),
	.B(B),
	.A_stb(A_stb),
    	.B_stb(B_stb),
	.result(Res),
	.result_ack(result_ack),
	.result_ready(ready)
);

 initial 
    begin
      forever
        #5 clk = !clk;
    end 

initial
  begin
    $monitor("Res_1_1=%b  \n Res_1_2=%b \n Res_1_3=%b",Res[1*FLOAT_SIZE-1:0*FLOAT_SIZE],Res[2*FLOAT_SIZE-1:1*FLOAT_SIZE],Res[3*FLOAT_SIZE-1:2*FLOAT_SIZE]);
    A = {16{one}};
    B = {16{one}};
    A_stb = 1'b1;
    B_stb = 1'b1;
    #15000;
    result_ack = 1'b1;
    A = 512'b01000000100010011001100110011010001111111100110011001100110011010011111011001100110011001100110100111110100110011001100110011010001111100100110011001100110011010100000011101001100110011001101001000000101110011001100110011010010000001010011001100110011001100100000011001001100110011001101001000000001000000000000000000000010000001001011001100110011001100100000000000110011001100110011001000000101010011001100110011010001111101100110011001100110011010100000000010011001100110011001100111111110000000000000000000000;
    B = 512'b01000000001000000000000000000000010000001101110011001100110011010100000000111001100110011001101001000000100011001100110011001101010000000111100110011001100110100100000010110011001100110011001101000001000111100110011001100110010000000101001100110011001100110100000011110110011001100110011001000000101000110011001100110011001111111010011001100110011001100011111111001100110011001100110101000000000001100110011001100110001111111111001100110011001100110011111111011001100110011001101000111111100011001100110011001101;
    A_stb = 1'b1;
    B_stb = 1'b1;
    #15000  $stop; 
  end 
  
endmodule